module multiplier_8x4bit(a,b,c);
input[7:0]a;
input[3:0]b;
output[11:0]c;
wire[11:0]w1,w2,w3,w4,w5,w6;
and(w1[0],a[0],b[0]);
and(w1[1],a[1],b[0]);
and(w1[2],a[2],b[0]);
and(w1[3],a[3],b[0]);
and(w1[4],a[4],b[0]);
and(w1[5],a[5],b[0]);
and(w1[6],a[6],b[0]);
and(w1[7],a[7],b[0]);
not(w1[8],1'b1);
not(w1[9],1'b1);
not(w1[10],1'b1);
not(w1[11],1'b1);
and(w2[1],a[0],b[1]);
and(w2[2],a[1],b[1]);
and(w2[3],a[2],b[1]);
and(w2[4],a[3],b[1]);
and(w2[5],a[4],b[1]);
and(w2[6],a[5],b[1]);
and(w2[7],a[6],b[1]);
and(w2[8],a[7],b[1]);
not(w2[0],1'b1);
not(w2[9],1'b1);
not(w2[10],1'b1);
not(w2[11],1'b1);
and(w3[2],a[0],b[2]);
and(w3[3],a[1],b[2]);
and(w3[4],a[2],b[2]);
and(w3[5],a[3],b[2]);
and(w3[6],a[4],b[2]);
and(w3[7],a[5],b[2]);
and(w3[8],a[6],b[2]);
and(w3[9],a[7],b[2]);
not(w3[0],1'b1);
not(w3[1],1'b1);
not(w3[10],1'b1);
not(w3[11],1'b1);
and(w4[3],a[0],b[3]);
and(w4[4],a[1],b[3]);
and(w4[5],a[2],b[3]);
and(w4[6],a[3],b[3]);
and(w4[7],a[4],b[3]);
and(w4[8],a[5],b[3]);
and(w4[9],a[6],b[3]);
and(w4[10],a[7],b[3]);
not(w4[0],1'b1);
not(w4[1],1'b1);
not(w4[2],1'b1);
not(w4[11],1'b1);
adder_12bit a1(w5,w1,w2);
adder_12bit a2(w6,w5,w3);
adder_12bit a3(c,w6,w4);
endmodule