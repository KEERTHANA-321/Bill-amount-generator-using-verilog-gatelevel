module rtshift(a,b,ed);
input [12:0]a;
input ed;
output [12:0]b;
wire[11:0]w;
and(w[0],a[2],a[2]);
and(b[0],ed,w[0]);
and(w[1],a[3],a[3]);
and(b[1],ed,w[1]);
and(w[2],a[4],a[4]);
and(b[2],ed,w[2]);
and(w[3],a[5],a[5]);
and(b[3],ed,w[3]);
and(w[4],a[6],a[6]);
and(b[4],ed,w[4]);
and(w[5],a[7],a[7]);
and(b[5],ed,w[5]);
and(w[6],a[8],a[8]);
and(b[6],ed,w[6]);
and(w[7],a[9],a[9]);
and(b[7],ed,w[7]);
and(w[8],a[10],a[10]);
and(b[8],ed,w[8]);
and(w[9],a[11],a[11]);
and(b[9],ed,w[9]);
and(w[10],a[12],a[12]);
and(b[10],ed,w[10]);
not(b[11],1'b1);
not(b[12],1'b1);
endmodule